

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity hardsigmoid is
  Port ( 
        data_in     : in std_logic_vector;
        data_out    : out std_logic_vector
  );
end hardsigmoid;

architecture Behavioral of hardsigmoid is

begin




end Behavioral;
